// arith_machine: execute a series of arithmetic instructions from an instruction cache
//
// except (output) - set to 1 when an unrecognized instruction is to be executed.
// clock  (input)  - the clock signal
// reset  (input)  - set to 1 to set all registers to zero, set to 0 for normal execution.

module arith_machine(except, clock, reset);
    output      except;
    input       clock, reset;
      
    wire [31:0] inst, rsData, rtData,B,imm32;  
    wire [31:0] PC,nextPC,out,out2;
    wire   overflow, zero, negative,overflow2, zero2, negative2;   
    wire [2:0] alu_op;
    wire       writeenable, rd_src, alu_src2;
    wire [4:0] rdNum;
    // DO NOT comment out or rename this module
    // or the test bench will break
    register #(32) PC_reg(PC, nextPC, clock, 1, reset);

    // DO NOT comment out or rename this module
    // or the test bench will break
    instruction_memory im(inst,PC[31:2]);

    // DO NOT comment out or rename this module
    // or the test bench will break
    regfile rf ( rsData, rtData,
                inst[25:21], inst[20:16], rdNum, out2, 
                writeenable, clock, reset);
    
    mips_decode mp(alu_op, writeenable, rd_src, alu_src2, except, inst[31:26], inst[5:0]);   
    /* add other modules */
    
    alu32 A1(nextPC, overflow, zero, negative, PC,32'h00000004, 3'b010);  
    
    mux2v mx1(B,rtData,imm32,alu_src2);  

    assign imm32 = {{16{inst[15]}}, inst[15:0]};

    mux2v #(5) mx0(rdNum, inst[15:11] ,inst[20:16],rd_src);


    alu32 A2(out2, overflow2, zero2, negative2, rsData, B , alu_op[2:0]);
endmodule // arith_machine
